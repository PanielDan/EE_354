//LFSR Code

module lfsr    (
out             ,  // Output of the counter
enable          ,  // Enable  for counter
clk             ,  // clock input
reset              // reset input
);

	output [7:0] out;

	input [7:0] data;
	input enable, clk, reset;
	reg [7:0] out;
	wire        linear_feedback;

	assign linear_feedback = !(out[7] ^ out[3]);

	always @(posedge clk)
	begin
		if (reset)
		out <= 8'b0 ;
		else if (enable) 
		begin
			out <= {out[6],out[5],
					out[4],out[3],
					out[2],out[1],
					out[0], linear_feedback};
		end 
	end
endmodule // End Of Module counter
